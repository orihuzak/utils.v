module utils

fn test_is_wsl() {
	assert is_wsl() == true
}
